
/* 
Full Adder Module for bit Addition 
Written by referencedesigner.com 
*/
`timescale 1ns / 100ps 
`include "shapeInt.v"

module tb_shapeInt; 
  // Declare inputs as regs and outputs as wires
  parameter N = 16;
  reg clock, reset;
  reg signed [N-1:0] data;
  wire signed [N-1:0] out;
  reg signed [N-1:0] Mpos=(1<<(N-1)) - 1;
  reg signed [N-1:0] Mneg=(1<<(N-1));
 
  shapeInt uut (
    .C(clock),
    .CLR(reset),
    .D(data),
    .Q(out)
  );
 

// Initialize all variables
initial 
  begin
   $display ( "time, ck, clr, data, out" );
   $monitor ( "%g, %b, %b, %d, %d" , $time, clock, reset, data, out);
   clock = 1; // initial value of clock
   reset = 0; // initial value of reset
   data = 0; // initial value of enable
   #5 reset = 1; // Assert the reset
   #10 reset = 0; // Deassert the reset
   #5 data = 0;
   #5 data =1024;
   #5 data =1013;
   #5 data =1003;
   #5 data =993;
   #5 data =983;
   #5 data =974;
   #5 data =964;
   #5 data =954;
   #5 data =945;
   #5 data =935;
   #5 data =926;
   #5 data =917;
   #5 data =908;
   #5 data =899;
   #5 data =890;
   #5 data =881;
   #5 data =872;
   #5 data =863;
   #5 data =855;
   #5 data =846;
   #5 data =838;
   #5 data =830;
   #5 data =821;
   #5 data =813;
   #5 data =805;
   #5 data =797;
   #5 data =789;
   #5 data =781;
   #5 data =773;
   #5 data =766;
   #5 data =758;
   #5 data =751;
   #5 data =743;
   #5 data =736;
   #5 data =728;
   #5 data =721;
   #5 data =714;
   #5 data =707;
   #5 data =700;
   #5 data =693;
   #5 data =686;
   #5 data =679;
   #5 data =672;
   #5 data =666;
   #5 data =659;
   #5 data =652;
   #5 data =646;
   #5 data =640;
   #5 data =633;
   #5 data =627;
   #5 data =621;
   #5 data =614;
   #5 data =608;
   #5 data =602;
   #5 data =596;
   #5 data =590;
   #5 data =584;
   #5 data =579;
   #5 data =573;
   #5 data =567;
   #5 data =561;
   #5 data =556;
   #5 data =550;
   #5 data =545;
   #5 data =539;
   #5 data =534;
   #5 data =529;
   #5 data =523;
   #5 data =518;
   #5 data =513;
   #5 data =508;
   #5 data =503;
   #5 data =498;
   #5 data =493;
   #5 data =488;
   #5 data =483;
   #5 data =478;
   #5 data =474;
   #5 data =469;
   #5 data =464;
   #5 data =460;
   #5 data =455;
   #5 data =451;
   #5 data =446;
   #5 data =442;
   #5 data =437;
   #5 data =433;
   #5 data =429;
   #5 data =424;
   #5 data =420;
   #5 data =416;
   #5 data =412;
   #5 data =408;
   #5 data =404;
   #5 data =400;
   #5 data =396;
   #5 data =392;
   #5 data =388;
   #5 data =384;
   #5 data =380;
   #5 data =376;
   #5 data =372;
   #5 data =369;
   #5 data =365;
   #5 data =361;
   #5 data =358;
   #5 data =354;
   #5 data =351;
   #5 data =347;
   #5 data =344;
   #5 data =340;
   #5 data =337;
   #5 data =334;
   #5 data =330;
   #5 data =327;
   #5 data =324;
   #5 data =321;
   #5 data =317;
   #5 data =314;
   #5 data =311;
   #5 data =308;
   #5 data =305;
   #5 data =302;
   #5 data =299;
   #5 data =296;
   #5 data =293;
   #5 data =290;
   #5 data =287;
   #5 data =284;
   #5 data =281;
   #5 data =279;
   #5 data =276;
   #5 data =273;
   #5 data =270;
   #5 data =268;
   #5 data =265;
   #5 data =262;
   #5 data =260;
   #5 data =257;
   #5 data =255;
   #5 data =252;
   #5 data =250;
   #5 data =247;
   #5 data =245;
   #5 data =242;
   #5 data =240;
   #5 data =237;
   #5 data =235;
   #5 data =233;
   #5 data =230;
   #5 data =228;
   #5 data =226;
   #5 data =223;
   #5 data =221;
   #5 data =219;
   #5 data =217;
   #5 data =215;
   #5 data =213;
   #5 data =210;
   #5 data =208;
   #5 data =206;
   #5 data =204;
   #5 data =202;
   #5 data =200;
   #5 data =198;
   #5 data =196;
   #5 data =194;
   #5 data =192;
   #5 data =190;
   #5 data =188;
   #5 data =187;
   #5 data =185;
   #5 data =183;
   #5 data =181;
   #5 data =179;
   #5 data =177;
   #5 data =176;
   #5 data =174;
   #5 data =172;
   #5 data =170;
   #5 data =169;
   #5 data =167;
   #5 data =165;
   #5 data =164;
   #5 data =162;
   #5 data =161;
   #5 data =159;
   #5 data =157;
   #5 data =156;
   #5 data =154;
   #5 data =153;
   #5 data =151;
   #5 data =150;
   #5 data =148;
   #5 data =147;
   #5 data =145;
   #5 data =144;
   #5 data =142;
   #5 data =141;
   #5 data =139;
   #5 data =138;
   #5 data =137;
   #5 data =135;
   #5 data =134;
   #5 data =133;
   #5 data =131;
   #5 data =130;
   #5 data =129;
   #5 data =127;
   #5 data =126;
   #5 data =125;
   #5 data =124;
   #5 data =122;
   #5 data =121;
   #5 data =120;
   #5 data =119;
   #5 data =118;
   #5 data =116;
   #5 data =115;
   #5 data =114;
   #5 data =113;
   #5 data =112;
   #5 data =111;
   #5 data =110;
   #5 data =109;
   #5 data =107;
   #5 data =106;
   #5 data =105;
   #5 data =104;
   #5 data =103;
   #5 data =102;
   #5 data =101;
   #5 data =100;
   #5 data =99;
   #5 data =98;
   #5 data =97;
   #5 data =96;
   #5 data =95;
   #5 data =94;
   #5 data =93;
   #5 data =92;
   #5 data =91;
   #5 data =91;
   #5 data =90;
   #5 data =89;
   #5 data =88;
   #5 data =87;
   #5 data =86;
   #5 data =85;
   #5 data =84;
   #5 data =84;
   #5 data =83;
   #5 data =82;
   #5 data =81;
   #5 data =80;
   #5 data =79;
   #5 data =79;
   #5 data =78;
   #5 data =77;
   #5 data =76;
   #5 data =76;
   #5 data =75;
   #5 data =74;
   #5 data =73;
   #5 data =73;
   #5 data =72;
   #5 data =71;
   #5 data =70;
   #5 data =70;
   #5 data =69;
   #5 data =68;
   #5 data =68;
   #5 data =67;
   #5 data =66;
   #5 data =66;
   #5 data =65;
   #5 data =64;
   #5 data =64;
   #5 data =63;
   #5 data =62;
   #5 data =62;
   #5 data =61;
   #5 data =61;
   #5 data =60;
   #5 data =59;
   #5 data =59;
   #5 data =58;
   #5 data =58;
   #5 data =57;
   #5 data =56;
   #5 data =56;
   #5 data =55;
   #5 data =55;
   #5 data =54;
   #5 data =54;
   #5 data =53;
   #5 data =53;
   #5 data =52;
   #5 data =52;
   #5 data =51;
   #5 data =50;
   #5 data =50;
   #5 data =49;
   #5 data =49;
   #5 data =48;
   #5 data =48;
   #5 data =48;
   #5 data =47;
   #5 data =47;
   #5 data =46;
   #5 data =46;
   #5 data =45;
   #5 data =45;
   #5 data =44;
   #5 data =44;
   #5 data =43;
   #5 data =43;
   #5 data =43;
   #5 data =42;
   #5 data =42;
   #5 data =41;
   #5 data =41;
   #5 data =40;
   #5 data =40;
   #5 data =40;
   #5 data =39;
   #5 data =39;
   #5 data =38;
   #5 data =38;
   #5 data =38;
   #5 data =37;
   #5 data =37;
   #5 data =37;
   #5 data =36;
   #5 data =36;
   #5 data =35;
   #5 data =35;
   #5 data =35;
   #5 data =34;
   #5 data =34;
   #5 data =34;
   #5 data =33;
   #5 data =33;
   #5 data =33;
   #5 data =32;
   #5 data =32;
   #5 data =32;
   #5 data =31;
   #5 data =31;
   #5 data =31;
   #5 data =30;
   #5 data =30;
   #5 data =30;
   #5 data =30;
   #5 data =29;
   #5 data =29;
   #5 data =29;
   #5 data =28;
   #5 data =28;
   #5 data =28;
   #5 data =27;
   #5 data =27;
   #5 data =27;
   #5 data =27;
   #5 data =26;
   #5 data =26;
   #5 data =26;
   #5 data =26;
   #5 data =25;
   #5 data =25;
   #5 data =25;
   #5 data =25;
   #5 data =24;
   #5 data =24;
   #5 data =24;
   #5 data =24;
   #5 data =23;
   #5 data =23;
   #5 data =23;
   #5 data =23;
   #5 data =22;
   #5 data =22;
   #5 data =22;
   #5 data =22;
   #5 data =22;
   #5 data =21;
   #5 data =21;
   #5 data =21;
   #5 data =21;
   #5 data =20;
   #5 data =20;
   #5 data =20;
   #5 data =20;
   #5 data =20;
   #5 data =19;
   #5 data =19;
   #5 data =19;
   #5 data =19;
   #5 data =19;
   #5 data =18;
   #5 data =18;
   #5 data =18;
   #5 data =18;
   #5 data =18;
   #5 data =18;
   #5 data =17;
   #5 data =17;
   #5 data =17;
   #5 data =17;
   #5 data =17;
   #5 data =16;
   #5 data =16;
   #5 data =16;
   #5 data =16;
   #5 data =16;
   #5 data =16;
   #5 data =15;
   #5 data =15;
   #5 data =15;
   #5 data =15;
   #5 data =15;
   #5 data =15;
   #5 data =15;
   #5 data =14;
   #5 data =14;
   #5 data =14;
   #5 data =14;
   #5 data =14;
   #5 data =14;
   #5 data =14;
   #5 data =13;
   #5 data =13;
   #5 data =13;
   #5 data =13;
   #5 data =13;
   #5 data =13;
   #5 data =13;
   #5 data =12;
   #5 data =12;
   #5 data =12;
   #5 data =12;
   #5 data =12;
   #5 data =12;
   #5 data =12;
   #5 data =12;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =11;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =10;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =9;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =8;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =7;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =6;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =5;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =4;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =3;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =2;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =1;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 data =0;
   #5 $finish;
  end

// Clock generator
always begin
#5 clock = ~clock; // Toggle clock every 5 ticks
end
 
endmodule
